module vect_mem_tb;


logic clk,we;
logic [31:0] a; 
logic [255:0]wd;
logic [255:0] rd;

vectmanager mem(clk,we,a,wd,rd);

initial begin
clk = 0;
# 10;
clk = 1;
we = 1;
a = 0;
wd = 256'b1111010101011111_0110111101101011_0100101010101000_0110111101101011_1111010101011111_0110111101101011_0100101010101000_0110111101101011_1111010101011111_0110111101101011_0100101010101000_0110111101101011_1111010101011111_0110111101101011_0100101010101000_0110111101101011;
#10;
clk = 0;
#10;
clk = 1;
we = 1;
a = 16;
wd = 256'b1111010101011111_0110111101101011_0100101010101000_0110111101101011_1111010101011111_0110111101101011_0100101010101000_0110111101101011_1111010101011111_0110111101101011_0100101010101000_0110111101101011_1111010101011111_0110111101101011_0100101010101000_0110111101101011;
#10;
clk = 0;
#10;
clk = 1;
we = 0;
a = 7;
#10;
end
endmodule